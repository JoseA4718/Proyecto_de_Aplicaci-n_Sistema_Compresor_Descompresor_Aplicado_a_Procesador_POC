module register_file(
	input [3:0] RS1,
	input [3:0] RS2,
	input [3:0] RS3,
	input [3:0] RD,
	input [31:0] WD,
	input wr_enable,
	input clk,
	input rst,
	
	output [31:0] RD1,
	output [31:0] RD2,
	output [31:0] RD3
	);
	
	logic [31:0] R0, R1, R2, R3, R4, R5, R6, R7, R8, R9, R10, R11, R12, R13, R14, R15;

	logic [31:0] RD1_temp, RD2_temp, RD3_temp;
	

	always @(*) begin
		
		case (RS1)
		
			// Reads register RS1
			4'd0: RD1_temp = R0; 	// register 0
			4'd1: RD1_temp = R1; 	// register 1
			4'd2: RD1_temp = R2; 	// register 2
			4'd3: RD1_temp = R3; 	// register 3
			4'd4: RD1_temp = R4; 	// register 4
			4'd5: RD1_temp = R5; 	// register 5
			4'd6: RD1_temp = R6; 	// register 6
			4'd7: RD1_temp = R7; 	// register 7
			4'd8: RD1_temp = R8; 	// register 8
			4'd9: RD1_temp = R9; 	// register 9
			4'd10: RD1_temp = R10; 	// register 10
			4'd11: RD1_temp = R11; 	// register 11
			4'd12: RD1_temp = R12; 	// register 12
			4'd13: RD1_temp = R13; 	// register 13
			4'd14: RD1_temp = R14; 	// register 14
			4'd15: RD1_temp = R15; 	// register 15
			default: RD1_temp = 0;
		
		endcase
		
		
		case (RS2)
		
			// Reads register RS2
			4'd0: RD2_temp = R0; // register 0
			4'd1: RD2_temp = R1; // register 1
			4'd2: RD2_temp = R2; // register 2
			4'd3: RD2_temp = R3; // register 3
			4'd4: RD2_temp = R4; // register 4
			4'd5: RD2_temp = R5; // register 5
			4'd6: RD2_temp = R6; // register 6
			4'd7: RD2_temp = R7; // register 7
			4'd8: RD2_temp = R8; // register 8
			4'd9: RD2_temp = R9; // register 9
			4'd10: RD2_temp = R10; // register 10
			4'd11: RD2_temp = R11; // register 11
			4'd12: RD2_temp = R12; // register 12
			4'd13: RD2_temp = R13; // register 13
			4'd14: RD2_temp = R14; // register 14
			4'd15: RD2_temp = R15; // register 15
			default: RD2_temp = 0;
		
		endcase
		
		
		case (RS3)
		
			// Reads register RS3
			4'd0: RD3_temp = R0; // register 0
			4'd1: RD3_temp = R1; // register 1
			4'd2: RD3_temp = R2; // register 2
			4'd3: RD3_temp = R3; // register 3
			4'd4: RD3_temp = R4; // register 4
			4'd5: RD3_temp = R5; // register 5
			4'd6: RD3_temp = R6; // register 6
			4'd7: RD3_temp = R7; // register 7
			4'd8: RD3_temp = R8; // register 8
			4'd9: RD3_temp = R9; // register 9
			4'd10: RD3_temp = R10; // register 10
			4'd11: RD3_temp = R11; // register 11
			4'd12: RD3_temp = R12; // register 12
			4'd13: RD3_temp = R13; // register 13
			4'd14: RD3_temp = R14; // register 14
			4'd15: RD3_temp = R15; // register 15
			default: RD3_temp = 0;
		
		endcase
		
	end
	
	always_ff @(posedge clk or posedge rst) begin
	
		if(rst)
		begin
			R0 = 32'd0;
			R1 = 32'd0;
			R2 = 32'd0;
			R3 = 32'd0;
			R4 = 32'd0;
			R5 = 32'd0;
			R6 = 32'd0;
			R7 = 32'd0;
			R8 = 32'd0;
			R9 = 32'd0;
			R10 = 32'd0;
			R11 = 32'd0;
			R12 = 32'd0;
			R13 = 32'd0;
			R14 = 32'd0;
			R15 = 32'd0;
		
		end
	
		else if (wr_enable)
		begin
		
			case (RD)
			
				// writes on A3 register
				4'd0: R0 = 31'd0; // register 0
				4'd1: R1 = WD; // register 1
				4'd2: R2 = WD; // register 2
				4'd3: R3 = WD; // register 3
				4'd4: R4 = WD; // register 4
				4'd5: R5 = WD; // register 5
				4'd6: R6 = WD; // register 6
				4'd7: R7 = WD; // register 7
				4'd8: R8 = WD; // register 8
				4'd9: R9 = WD; // register 9
				4'd10: R10 = WD; // register 10
				4'd11: R11 = WD; // register 11
				4'd12: R12 = WD; // register 12
				4'd13: R13 = WD; // register 13
				4'd14: R14 = WD; // register 14
				4'd15: R15 = WD;
			
			endcase
		
		end
		
		
		
	end
		
		
	// output logic
	assign RD1 = RD1_temp;
	assign RD2 = RD2_temp;
	assign RD3 = RD3_temp;

	
endmodule